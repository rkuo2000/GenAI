* RC Low-Pass Filter
V1 in 0 AC 1 SIN(0 1 1k)
R1 in out 1k
C1 out 0 1uF

.AC DEC 10 10 100k

.control
set gnuplot_terminal="png"
run
gnuplot gp v(out) v(in)
.endc
.END
